`timescale 1ns / 1ps

module ALUController (
    //Inputs
    input logic [1:0] ALUOp,  // 2-bit opcode field from the Controller--00: LW/SW/AUIPC; 01:Branch; 10: Rtype/Itype; 11:JAL/LUI
    input logic [6:0] Funct7,  // bits 25 to 31 of the instruction
    input logic [2:0] Funct3,  // bits 12 to 14 of the instruction

    //Output
    output logic [3:0] Operation  // operation selection for ALU
);

  assign Operation[0] = 
                              (ALUOp == 2'b00) ||                                                    // load, store
                              ((ALUOp == 2'b10) && (Funct3 == 3'b110)) ||                            // or, ori
                              ((ALUOp == 2'b10) && (Funct3 == 3'b000) && (Funct7 == 7'b0000000)) ||  // add
                              ((ALUOp == 2'b10) && (Funct3 == 3'b000) && (Funct7 != 7'b0100000)) ||  // addi
                              ((ALUOp == 2'b10) && (Funct3 == 3'b101) && (Funct7 == 7'b0000000)) ||  // srl, srli
                              ((ALUOp == 2'b10) && (Funct3 == 3'b001) && (Funct7 == 7'b0000000)) ||  // sll, slli
                              ((ALUOp == 2'b01) && (Funct3 == 3'b001)) ||                            // bne
                              ((ALUOp == 2'b01) && (Funct3 == 3'b100)) ||                            // blt
                              ((ALUOp == 2'b01) && (Funct3 == 3'b101)) ||                            // bge
                              ((ALUOp == 2'b01) && (Funct3 == 3'b111)) ||                            // bgeu
                              (ALUOp == 2'b11);                                                      // lui

  assign Operation[1] = 
                              (ALUOp == 2'b00) ||                                                    // LOAD, STORE
                              ((ALUOp == 2'b10) && (Funct3 == 3'b100)) ||                            // XOR, XORI
                              ((ALUOp == 2'b10) && (Funct3 == 3'b000) && (Funct7 == 7'b0000000)) ||  // ADD
                              ((ALUOp == 2'b10) && (Funct3 == 3'b000) && (Funct7 != 7'b0100000)) ||  // ADDI
                              ((ALUOp == 2'b10) && (Funct3 == 3'b101) && (Funct7 == 7'b0100000)) ||  // SRA, SRAI
                              ((ALUOp == 2'b10) && (Funct3 == 3'b001) && (Funct7 == 7'b0000000)) ||  // SLL, SLLI
                              ((ALUOp == 2'b10) && (Funct3 == 3'b010)) ||                            // SLT, SLTI
                              ((ALUOp == 2'b01) && (Funct3 == 3'b101)) ||                            // BGE
                              ((ALUOp == 2'b01) && (Funct3 == 3'b110)) ||                            // BLTU
                              ((ALUOp == 2'b10) && (Funct3 == 3'b011)) ||                            // SLTU, SLTIU
                              ((ALUOp == 2'b01) && (Funct3 == 3'b111));                              // BGEU



  assign Operation[2] = 
                              ((ALUOp == 2'b10) && (Funct3 == 3'b000) && (Funct7 == 7'b0100000)) ||  // SUB
                              ((ALUOp == 2'b10) && (Funct3 == 3'b101) && (Funct7 == 7'b0000000)) ||  // SRL, SRLI
                              ((ALUOp == 2'b10) && (Funct3 == 3'b101) && (Funct7 == 7'b0100000)) ||  // SRA, SRAI
                              ((ALUOp == 2'b10) && (Funct3 == 3'b001) && (Funct7 == 7'b0000000)) ||  // SLL, SLLI
                              ((ALUOp == 2'b11) && (Funct3 == 3'b000)) ||                            // JALR
                              ((ALUOp == 2'b01) && (Funct3 == 3'b110)) ||                            // BLTU
                              ((ALUOp == 2'b10) && (Funct3 == 3'b011)) ||                            // SLTU, SLTIU
                              ((ALUOp == 2'b01) && (Funct3 == 3'b111)) ||                            // BGEU
                              (ALUOp == 2'b11);                                                      // LUI



  assign Operation[3] = 
                              ((ALUOp == 2'b01) && (Funct3 == 3'b000)) ||                            // BEQ
                              ((ALUOp == 2'b01) && (Funct3 == 3'b001)) ||                            // BNE
                              ((ALUOp == 2'b01) && (Funct3 == 3'b100)) ||                            // BLT
                              ((ALUOp == 2'b01) && (Funct3 == 3'b101)) ||                            // BGE
                              ((ALUOp == 2'b10) && (Funct3 == 3'b010)) ||                            // SLT, SLTI
                              ((ALUOp == 2'b11) && (Funct3 == 3'b000)) ||                            // JALR
                              ((ALUOp == 2'b01) && (Funct3 == 3'b110)) ||                            // BLTU
                              ((ALUOp == 2'b10) && (Funct3 == 3'b011)) ||                            // SLTU, SLTIU
                              ((ALUOp == 2'b01) && (Funct3 == 3'b111)) ||                            // BGEU
                              (ALUOp == 2'b11);                                                      // LUI
endmodule
